/*
 Data Encryption Standard (S-DES)
 64-bit 16-round block cipher encryption and decryption algorithm 
 using 56-bit key (64-bit key with Parity).
 */

module GenerateKeys (Key, SubKey1, SubKey2, SubKey3, SubKey4,
		     SubKey5, SubKey6, SubKey7, SubKey8,
		     SubKey9, SubKey10, SubKey11, SubKey12,
		     SubKey13, SubKey14, SubKey15, SubKey16);
   
   // Generate SubKeys
   input logic [63:0]  Key;
   output logic [47:0] SubKey1;
   output logic [47:0] SubKey2;
   output logic [47:0] SubKey3;
   output logic [47:0] SubKey4;
   output logic [47:0] SubKey5;
   output logic [47:0] SubKey6;
   output logic [47:0] SubKey7;
   output logic [47:0] SubKey8;
   output logic [47:0] SubKey9;
   output logic [47:0] SubKey10;
   output logic [47:0] SubKey11;
   output logic [47:0] SubKey12;
   output logic [47:0] SubKey13;
   output logic [47:0] SubKey14;
   output logic [47:0] SubKey15;
   output logic [47:0] SubKey16;
   
   //IP
   logic [27:0] left_block, right_block;
   logic [27:0] lb1, lb2, lb3, lb4, lb5, lb6, lb7, lb8, lb9, lb10, lb11, lb12, lb13, lb14, lb15, lb16;
   logic [27:0] rb1, rb2, rb3, rb4, rb5, rb6, rb7, rb8, rb9. rb10, rb11, rb12, rb13, rb14, rb15, rb16;

<<<<<<< HEAD
   PC1 mod1(Key, left_block, right_block); //first scrambled then cut in half

   assign lb1 = {left_block[26:0], left_block[27]}; //shift left and right block by 1
   assign rb1 = {right_block[26:0], right_block[27]}; 

   PC2 mod2(lb1, rb1, subkey1); //scrambled combined left/right blocks to get subkey1

   assign lb2 = {lb1[26:0], lb1[27]}; //shift new left/right blocks by 1
   assign rb2 = {rb1[26:0], rb1[27]};

   PC2 mod3(lb2, rb2, subkey2); //scrambled combined new left/right blocks to get subkey2

   assign lb3 = {lb2[25:0], lb2[27:26]}; //shift new left/right blocks by 2
   assign rb3 = {rb2[25:0], rb2[27:26]};
   
   PC2 mod4(lb3, rb3, subkey3); //scrambled combined new left/right blocks to get subkey3
   
   assign lb4 = {lb3[25:0], lb3[27:26]}; //shift new left/right blocks by 2
   assign rb4 = {rb3[25:0], rb3[27:26]};
   
   PC2 mod5(lb4, rb4, subkey4); //scrambled combined new left/right blocks to get subkey4
   
   assign lb5 = {lb4[25:0], lb4[27:26]}; //shift new left/right blocks by 2
   assign rb5 = {rb4[25:0], rb4[27:26]};
   
   PC2 mod6(lb5, rb5, subkey5); //scrambled combined new left/right blocks to get subkey5
   
   assign lb6 = {lb5[25:0], lb5[27:26]}; //shift new left/right blocks by 2
   assign rb6 = {rb5[25:0], rb5[27:26]};
   
   PC2 mod7(lb6, rb6, subkey6); //scrambled combined new left/right blocks to get subkey6
   
   assign lb7 = {lb6[25:0], lb6[27:26]}; //shift new left/right blocks by 2
   assign rb7 = {rb6[25:0], rb6[27:26]};
   
   PC2 mod8(lb7, rb7, subkey7); //scrambled combined new left/right blocks to get subkey7
   
   assign lb8 = {lb7[25:0], lb7[27:26]}; //shift new left/right blocks by 2
   assign rb8 = {rb7[25:0], rb7[27:26]};

   PC2 mod9(lb8, rb8, subkey8); //scrambled combined new left/right blocks to get subkey8
   
   assign lb9 = {lb8[26:0], lb8[27]}; //shift new left/right blocks by 1
   assign rb9 = {rb8[26:0], rb8[27]};

   PC2 mod10(lb9, rb9, subkey9); //scrambled combined new left/right blocks to get subkey9
   
   assign lb10 = {lb9[25:0], lb9[27:26]}; //shift new left/right blocks by 2
   assign rb10 = {rb9[25:0], rb9[27:26]}; 
   
   PC2 mod11(lb10, rb10, subkey10); //scrambled combined new left/right blocks to get subkey10
   
   assign lb11 = {lb10[25:0], lb10[27:26]}; //shift new left/right blocks by 2
   assign rb11 = {rb10[25:0], rb10[27:26]};
   
   PC2 mod12(lb11, rb11, subkey11); //scrambled combined new left/right blocks to get subkey11
   
   assign lb12 = {lb11[25:0], lb11[27:26]}; //shift new left/right blocks by 2
   assign rb12 = {rb11[25:0], rb11[27:26]};
   
   PC2 mod13(lb12, rb12, subkey12); //scrambled combined new left/right blocks to get subkey12
   
   assign lb13 = {lb12[25:0], lb12[27:26]}; //shift new left/right blocks by 2
   assign rb13 = {rb12[25:0], rb12[27:26]};
   
   PC2 mod14(lb13, rb13, subkey13); //scrambled combined new left/right blocks to get subkey13
   
   assign lb14 = {lb13[25:0], lb13[27:26]}; //shift new left/right blocks by 2
   assign rb14 = {rb13[25:0], rb13[27:26]};
   
   PC2 mod15(lb14, rb14, subkey14); //scrambled combined new left/right blocks to get subkey14
   
   assign lb15 = {lb14[25:0], lb14[27:26]}; //shift new left/right blocks by 2
   assign rb15 = {rb14[25:0], rb14[27:26]};

   PC2 mod16(lb15, rb15, subkey15); //scrambled combined new left/right blocks to get subkey15
   
   assign rb16 = {rb15[26:0], rb15[27]}; //shift new left/right blocks by 1
   assign lb16 = {lb15[26:0], lb15[27]};

   PC2 mod17(lb16, rb16, subkey16);
=======
	//pc1 v1
   logic [27:0] left_block, right_block;
   logic [27:0] lb1, rb1;
   PC1 mod1(Key, left_block, right_block);
   assign lb1 = {left_block[54:28], left_block[55]};
   assign rb1 = {right_block[26:0], right_block[27]};
    //pc1 v2
   logic [27:0] lb2, rb2;
   PC2 mod2(lb1, rb1, subkey1);
   assign lb2 = {lb1[54:28], lb1[55]};
   assign rb2 = {rb1[26:0], rb1[27]};

    //pc1 v3
   logic [27:0] lb3, rb3;
   PC2 mod3(lb2, rb2, subkey2);
   assign lb3 = {lb2[53:28], lb2[55:54]};
   assign rb3 = {rb2[25:0], rb2[27:26]};
    //pc1 v4
   logic [27:0] lb4, rb4;
   PC2 mod4(lb3, rb3, subkey3);
   assign lb4 = {lb3[53:28], lb3[55:54]};
   assign rb4 = {rb3[25:0], rb3[27:26]};
    //pc1 v5
   logic [27:0] lb5, rb5;
   PC2 mod2(lb4, rb4, subkey4);
   assign lb5 = {lb4[53:28], lb4[55:54]};
   assign rb5 = {rb4[25:0], rb4[27:26]};
    //pc1 v6
   logic [27:0] lb6, rb6;
   PC2 mod2(lb5, rb5, subkey5);
   assign lb6 = {lb5[53:28], lb5[55:54]};
   assign rb6 = {rb5[25:0], rb5[27:26]};
    //pc1 v7
   logic [27:0] lb7, rb7;
   PC2 mod2(lb6, rb6, subkey6);
   assign lb7 = {lb6[53:28], lb6[55:54]};
   assign rb7 = {rb6[25:0], rb6[27:26]};
    //pc1 v8
   logic [27:0] lb8, rb8;
   PC2 mod2(lb7, rb7, subkey7);
   assign lb8 = {lb7[53:28], lb7[55:54]};
   assign rb8 = {rb7[25:0], rb7[27:26]};

    //pc1 v9
   logic [27:0] lb9, rb9;
   PC2 mod2(lb8, rb8, subkey8);
   assign lb9 = {lb8[54:28], lb8[55]};
   assign rb9 = {rb8[26:0], rb8[27]};

    //pc1 v10
   logic [27:0] lb10, rb10;
   PC2 mod2(lb9, rb9, subkey9);
   assign lb10 = {lb9[53:28], lb9[55:54]};
   assign rb10 = {rb9[26:0], rb9[27:26]}; 
    //pc1 v11
   logic [27:0] lb11, rb11;
   PC2 mod2(lb10, rb10, subkey10);
   assign lb11 = {lb10[53:28], lb10[55:54]};
   assign rb11 = {rb10[25:0], rb10[27:26]};
    //pc1 v12
   logic [27:0] lb12, rb12;
   PC2 mod2(lb11, rb11, subkey11);
   assign lb12 = {lb11[53:28], lb11[55:54]};
   assign rb12 = {rb11[25:0], rb11[27:26]};
    //pc1 v13
   logic [27:0] lb13, rb13;
   PC2 mod2(lb12, rb12, subkey12);
   assign lb13 = {lb12[53:28], lb12[55:54]};
   assign rb13 = {rb12[25:0], rb12[27:26]};
    //pc1 v14
   logic [27:0] lb14, rb14;
   PC2 mod2(lb13, rb13, subkey13);
   assign lb14 = {lb13[53:28], lb13[55:54]};
   assign rb14 = {rb13[25:0], rb13[27:26]};
    //pc1 v15
   logic [27:0] lb15, rb15;
   PC2 mod2(lb14, rb14, subkey14);
   assign lb15 = {lb14[53:28], lb14[55:54]};
   assign rb15 = {rb14[25:0], rb14[27:26]};

    //pc1 v16
   logic [27:0] lb16, rb16;
   PC2 mod2(lb15, rb15, subkey15);
   assign lb16 = {lb15[54:28], lb15[55]};
   assign rb16 = {rb15[26:0], rb15[27]};
>>>>>>> 2cb05479a716221d24a2dce71af84162bc87bae0

endmodule // GenerateKeys

module PC1 (key, left_block, right_block);

   input logic [63:0]  key;
   output logic [27:0] left_block;
   output logic [27:0] right_block;

   logic [55:0] out_block;

//left
   assign out_block[55] = key[64-57];
   assign out_block[54] = key[64-49];
   assign out_block[53] = key[64-41];
   assign out_block[52] = key[64-33];
   assign out_block[51] = key[64-25];
   assign out_block[50] = key[64-17];
   assign out_block[49] = key[64-9];
   assign out_block[48] = key[64-1];
   assign out_block[47] = key[64-58];
   assign out_block[46] = key[64-50];   
   assign out_block[45] = key[64-42];   
   assign out_block[44] = key[64-34];
   assign out_block[43] = key[64-26];
   assign out_block[42] = key[64-18];
   assign out_block[41] = key[64-10];
   assign out_block[40] = key[64-2];
   assign out_block[39] = key[64-59];
   assign out_block[38] = key[64-51];
   assign out_block[37] = key[64-43];
   assign out_block[36] = key[64-35];   
   assign out_block[35] = key[64-27];
   assign out_block[34] = key[64-19];   
   assign out_block[33] = key[64-11];
   assign out_block[32] = key[64-3];
   assign out_block[31] = key[64-60];
   assign out_block[30] = key[64-52];
   assign out_block[29] = key[64-44];
   assign out_block[28] = key[64-36];


   //right
   assign out_block[27] = key[64-63];
   assign out_block[26] = key[64-55];   
   assign out_block[25] = key[64-47];
   assign out_block[24] = key[64-39];   
   assign out_block[23] = key[64-31];
   assign out_block[22] = key[64-23];
   assign out_block[21] = key[64-15];
   assign out_block[20] = key[64-7];
   assign out_block[19] = key[64-62];
   assign out_block[18] = key[64-54];
   assign out_block[17] = key[64-46];   
   assign out_block[16] = key[64-38];   
   assign out_block[15] = key[64-30];
   assign out_block[14] = key[64-22];   
   assign out_block[13] = key[64-14];
   assign out_block[12] = key[64-6];
   assign out_block[11] = key[64-61];
   assign out_block[10] = key[64-53];
   assign out_block[9] = key[64-45];
   assign out_block[8] = key[64-37];
   assign out_block[7] = key[64-29];
   assign out_block[6] = key[64-21];   
   assign out_block[5] = key[64-13];
   assign out_block[4] = key[64-5];   
   assign out_block[3] = key[64-28];
   assign out_block[2] = key[64-20];
   assign out_block[1] = key[64-12];
   assign out_block[0] = key[64-4];
   
endmodule // PC1

module PC2 (left_block, right_block, subkey);

   input logic [27:0] left_block;
   input logic [27:0] right_block;
   output logic [47:0] subkey;
   
   logic [47:0] combined;

   assign combined = {left_block, right};
   
   assign subkey[47] = combined[56-14];
   assign subkey[46] = combined[56-17];
   assign subkey[45] = combined[56-11];
   assign subkey[44] = combined[56-24];   
   assign subkey[43] = combined[56-1];
   assign subkey[42] = combined[56-5];   
   assign subkey[41] = combined[56-3];
   assign subkey[40] = combined[56-28];
   assign subkey[39] = combined[56-15];
   assign subkey[38] = combined[56-6];
   assign subkey[37] = combined[56-21];
   assign subkey[36] = combined[56-10];
   assign subkey[35] = combined[56-23];
   assign subkey[34] = combined[56-19];   
   assign subkey[33] = combined[56-12];
   assign subkey[32] = combined[56-4];   
   assign subkey[31] = combined[56-26];
   assign subkey[30] = combined[56-8];
   assign subkey[29] = combined[56-16];
   assign subkey[28] = combined[56-7];
   assign subkey[27] = combined[56-27];
   assign subkey[26] = combined[56-20];
   assign subkey[25] = combined[56-13];   
   assign subkey[24] = combined[56-2];   
   assign subkey[23] = combined[56-41];
   assign subkey[22] = combined[56-52];   
   assign subkey[21] = combined[56-31];
   assign subkey[20] = combined[56-37];
   assign subkey[19] = combined[56-47];
   assign subkey[18] = combined[56-55];
   assign subkey[17] = combined[56-30];
   assign subkey[16] = combined[56-40];
   assign subkey[15] = combined[56-51];
   assign subkey[14] = combined[56-45];   
   assign subkey[13] = combined[56-33];
   assign subkey[12] = combined[56-48];   
   assign subkey[11] = combined[56-44];
   assign subkey[10] = combined[56-49];
   assign subkey[9] = combined[56-39];
   assign subkey[8] = combined[56-56];
   assign subkey[7] = combined[56-34];
   assign subkey[6] = combined[56-53];
   assign subkey[5] = combined[56-46];
   assign subkey[4] = combined[56-42];   
   assign subkey[3] = combined[56-50];
   assign subkey[2] = combined[56-36];    
   assign subkey[1] = combined[56-29];
   assign subkey[0] = combined[56-32];

endmodule // PC2

// Straight Function
module SF (inp_block, out_block);

   input logic [31:0] inp_block;
   output logic [31:0] out_block;

   assign out_block=[31] = inp_block[32-16];
   assign out_block=[30] = inp_block[32-7];
   assign out_block=[29] = inp_block[32-20];
   assign out_block=[28] = inp_block[32-21];
   assign out_block=[27] = inp_block[32-29];
   assign out_block=[26] = inp_block[32-12];
   assign out_block=[25] = inp_block[32-28];
   assign out_block=[24] = inp_block[32-17];
   assign out_block=[23] = inp_block[32-1];
   assign out_block=[22] = inp_block[32-15];
   assign out_block=[21] = inp_block[32-23];
   assign out_block=[20] = inp_block[32-26];
   assign out_block=[19] = inp_block[32-5];
   assign out_block=[18] = inp_block[32-18];
   assign out_block=[17] = inp_block[32-31];
   assign out_block=[16] = inp_block[32-10];
   assign out_block=[15] = inp_block[32-2];
   assign out_block=[14] = inp_block[32-8];
   assign out_block=[13] = inp_block[32-24];
   assign out_block=[12] = inp_block[32-14];
   assign out_block=[11] = inp_block[32-23];
   assign out_block=[10] = inp_block[32-27];
   assign out_block=[9] = inp_block[32-3];
   assign out_block=[8] = inp_block[32-9];
   assign out_block=[7] = inp_block[32-19];
   assign out_block=[6] = inp_block[32-13];
   assign out_block=[5] = inp_block[32-30];
   assign out_block=[4] = inp_block[32-6];
   assign out_block=[3] = inp_block[32-22];
   assign out_block=[2] = inp_block[32-11];
   assign out_block=[1] = inp_block[32-4];
   assign out_block=[0] = inp_block[32-25];

endmodule // SF

// Expansion Function
module EF (inp_block, out_block);

   input logic [31:0] inp_block;
   output logic [47:0] out_block;

   assign out_block=[46] = inp_block[32-32];
   assign out_block=[45] = inp_block[32-1];
   assign out_block=[44] = inp_block[32-2];
   assign out_block=[47] = inp_block[32-3];
   assign out_block=[43] = inp_block[32-4];
   assign out_block=[42] = inp_block[32-5];
   assign out_block=[41] = inp_block[32-4];
   assign out_block=[40] = inp_block[32-5];
   assign out_block=[39] = inp_block[32-6];
   assign out_block=[38] = inp_block[32-7];
   assign out_block=[37] = inp_block[32-8];
   assign out_block=[36] = inp_block[32-9];
   assign out_block=[35] = inp_block[32-8];
   assign out_block=[34] = inp_block[32-9];
   assign out_block=[33] = inp_block[32-10];
   assign out_block=[32] = inp_block[32-11];
   assign out_block=[31] = inp_block[32-12];
   assign out_block=[30] = inp_block[32-13];
   assign out_block=[29] = inp_block[32-12];
   assign out_block=[28] = inp_block[32-13];
   assign out_block=[27] = inp_block[32-14];
   assign out_block=[26] = inp_block[32-15];
   assign out_block=[25] = inp_block[32-16];
   assign out_block=[24] = inp_block[32-17];
   assign out_block=[23] = inp_block[32-16];
   assign out_block=[22] = inp_block[32-17];
   assign out_block=[21] = inp_block[32-18];
   assign out_block=[20] = inp_block[32-19];
   assign out_block=[19] = inp_block[32-20];
   assign out_block=[18] = inp_block[32-21];
   assign out_block=[17] = inp_block[32-20];
   assign out_block=[16] = inp_block[32-21];
   assign out_block=[15] = inp_block[32-22];
   assign out_block=[14] = inp_block[32-23];
   assign out_block=[13] = inp_block[32-24];
   assign out_block=[12] = inp_block[32-25];
   assign out_block=[11] = inp_block[32-24];
   assign out_block=[10] = inp_block[32-25];
   assign out_block=[9] = inp_block[32-26];
   assign out_block=[8] = inp_block[32-27];
   assign out_block=[7] = inp_block[32-28];
   assign out_block=[6] = inp_block[32-29];
   assign out_block=[5] = inp_block[32-28];
   assign out_block=[4] = inp_block[32-29];
   assign out_block=[3] = inp_block[32-30];
   assign out_block=[2] = inp_block[32-31];
   assign out_block=[1] = inp_block[32-32];
   assign out_block=[0] = inp_block[32-1];

endmodule // EF

module feistel (inp_block, subkey, out_block);

   input logic [31:0]  inp_block;
   input logic [47:0]  subkey;
   output logic [31:0] out_block;

<<<<<<< HEAD
   logic [47:0] e_inp; //expanded right block 1 from round
   logic [47:0] xe_inp; //XORed e_inp
   logic [31:0] bxe_inp; //boxed xe_inp

   EF feist(inp_block, e_inp); //scrambled
   
   assign xe_inp = e_inp ^ subkey;

   S8_Box s8(xe_inp[5:0], bxe_inp[3:0]);
   S7_Box s7(xe_inp[11:6], bxe_inp[7:4]);
   S6_Box s6(xe_inp[17:12], bxe_inp[11:8]);
   S5_Box s5(xe_inp[23:18], bxe_inp[15:12]);
   S4_Box s4(xe_inp[29:24], bxe_inp[19:16]);
   S3_Box s3(xe_inp[35:30], bxe_inp[23:20]);
   S2_Box s2(xe_inp[41:36], bxe_inp[27:24]);
   S1_Box s1(xe_inp[47:42], bxe_inp[31:28]);

   SF straight(bxe_inp, out_block); //scrambled
   
=======
   logic [47:0] e_inp; //expanded inp_block
   logic [47:0] xe_inp; //XORed e_inp
   logic [32:0] f_inp; //straight xe_inp

   EF feist(inp_block, e_inp);
   
   assign xe_inp = e_inp ^ subkey;

   S8_Box s8(xe_inp[5:0],f_inp[3:0]);
   S7_Box s7(xe_inp[11:6],f_inp[7:4]);
   S6_Box s6(xe_inp[17:12],f_inp[11:8]);
   S5_Box s5(xe_inp[23:18],f_inp[15:12]);
   S4_Box s4(xe_inp[29:24],f_inp[19:16]);
   S3_Box s3(xe_inp[35:30],f_inp[23:20]);
   S2_Box s2(xe_inp[41:36],f_inp[27:24]);
   S1_Box s1(xe_inp[47:42],f_inp[31:28]);

   SF straight(f_inp, xe_inp);
   

>>>>>>> 2cb05479a716221d24a2dce71af84162bc87bae0
endmodule // Feistel

// DES block round
module round (inp_block, subkey, out_block);

   input logic  [63:0]  inp_block;
   input logic  [47:0]  subkey;
<<<<<<< HEAD
   output logic [63:0]  out_block;

   logic [31:0] left_block1, right_block1;
   logic [31:0] left_block2, right_block2;
   logic [31:0] feisteled_block;

   assign left_block1 = inp_block[63:32];
   assign right_block1 = inp_block[31:0];

   feistel fb(rightblock1, subkey, feisteled_block);

   assign left_block2 = right_block1;
   assign right_block2 = feisteled_block ^ left_block1;
   assign out_block = {left_block2, right_block2};
=======
   output logic [63:0] out_block;
>>>>>>> 2cb05479a716221d24a2dce71af84162bc87bae0

   logic [31:0] left_block1, right_block1;
   logic [31:0] left_block2, right_block2;
   logic [31:0] feisteled_block;

   assign left_block1 = inp_block[63:32];
   assign right_block1 = inp_block[31:0];

   feistel fb(rightblock1, subkey, feisteled_block);

   assign left_block2 = right_block1;
   assign right_block2 = feisteled_block ^ left_block;
   assign out_block = {left_block2, right_block2};

endmodule // round1

// Initial Permutation
module IP (inp_block, out_block);

   input logic [63:0]  inp_block;
   output logic [63:0] out_block;

   assign out_block[63] = inp_block[64-58];
   assign out_block[62] = inp_block[64-50];
   assign out_block[61] = inp_block[64-42];
   assign out_block[60] = inp_block[64-34];
   assign out_block[59] = inp_block[64-26];
   assign out_block[58] = inp_block[64-18];
   assign out_block[57] = inp_block[64-10];
   assign out_block[56] = inp_block[64-2];
   assign out_block[55] = inp_block[64-60];
   assign out_block[54] = inp_block[64-52];   
   assign out_block[53] = inp_block[64-44];   
   assign out_block[52] = inp_block[64-36];
   assign out_block[51] = inp_block[64-28];
   assign out_block[50] = inp_block[64-20];
   assign out_block[49] = inp_block[64-12];
   assign out_block[48] = inp_block[64-4];
   assign out_block[47] = inp_block[64-62];
   assign out_block[46] = inp_block[64-54];
   assign out_block[45] = inp_block[64-46];
   assign out_block[44] = inp_block[64-38];   
   assign out_block[43] = inp_block[64-30];
   assign out_block[42] = inp_block[64-22];   
   assign out_block[41] = inp_block[64-14];
   assign out_block[40] = inp_block[64-6];
   assign out_block[39] = inp_block[64-64];
   assign out_block[38] = inp_block[64-56];
   assign out_block[37] = inp_block[64-48];
   assign out_block[36] = inp_block[64-40];
   assign out_block[35] = inp_block[64-32];
   assign out_block[34] = inp_block[64-24];   
   assign out_block[33] = inp_block[64-16];
   assign out_block[32] = inp_block[64-8];   
   assign out_block[31] = inp_block[64-57];
   assign out_block[30] = inp_block[64-49];
   assign out_block[29] = inp_block[64-41];
   assign out_block[28] = inp_block[64-33];
   assign out_block[27] = inp_block[64-25];
   assign out_block[26] = inp_block[64-17];
   assign out_block[25] = inp_block[64-9];   
   assign out_block[24] = inp_block[64-1];   
   assign out_block[23] = inp_block[64-59];
   assign out_block[22] = inp_block[64-51];   
   assign out_block[21] = inp_block[64-43];
   assign out_block[20] = inp_block[64-35];
   assign out_block[19] = inp_block[64-27];
   assign out_block[18] = inp_block[64-19];
   assign out_block[17] = inp_block[64-11];
   assign out_block[16] = inp_block[64-3];
   assign out_block[15] = inp_block[64-61];
   assign out_block[14] = inp_block[64-53];   
   assign out_block[13] = inp_block[64-45];
   assign out_block[12] = inp_block[64-37];   
   assign out_block[11] = inp_block[64-29];
   assign out_block[10] = inp_block[64-21];
   assign out_block[9] = inp_block[64-13];
   assign out_block[8] = inp_block[64-5];
   assign out_block[7] = inp_block[64-63];
   assign out_block[6] = inp_block[64-55];
   assign out_block[5] = inp_block[64-47];
   assign out_block[4] = inp_block[64-39];   
   assign out_block[3] = inp_block[64-31];
   assign out_block[2] = inp_block[64-23];    
   assign out_block[1] = inp_block[64-15];
   assign out_block[0] = inp_block[64-7];   

endmodule // IP

// Final Permutation
module FP (inp_block, out_block);

   input logic [63:0]  inp_block;
   output logic [63:0] out_block;

   assign out_block[63] = inp_block[64-40];
   assign out_block[62] = inp_block[64-8];
   assign out_block[61] = inp_block[64-48];
   assign out_block[60] = inp_block[64-16];
   assign out_block[59] = inp_block[64-56];
   assign out_block[58] = inp_block[64-24];
   assign out_block[57] = inp_block[64-64];
   assign out_block[56] = inp_block[64-32];   
   assign out_block[55] = inp_block[64-39];
   assign out_block[54] = inp_block[64-7];   
   assign out_block[53] = inp_block[64-47];   
   assign out_block[52] = inp_block[64-15];
   assign out_block[51] = inp_block[64-55];
   assign out_block[50] = inp_block[64-23];
   assign out_block[49] = inp_block[64-63];
   assign out_block[48] = inp_block[64-31];   
   assign out_block[47] = inp_block[64-38];
   assign out_block[46] = inp_block[64-6];
   assign out_block[45] = inp_block[64-46];
   assign out_block[44] = inp_block[64-14];   
   assign out_block[43] = inp_block[64-54];
   assign out_block[42] = inp_block[64-22];   
   assign out_block[41] = inp_block[64-62];
   assign out_block[40] = inp_block[64-30];   
   assign out_block[39] = inp_block[64-37];
   assign out_block[38] = inp_block[64-5];
   assign out_block[37] = inp_block[64-45];
   assign out_block[36] = inp_block[64-13];
   assign out_block[35] = inp_block[64-53];
   assign out_block[34] = inp_block[64-21];   
   assign out_block[33] = inp_block[64-61];
   assign out_block[32] = inp_block[64-29];   
   assign out_block[31] = inp_block[64-36];
   assign out_block[30] = inp_block[64-4];
   assign out_block[29] = inp_block[64-44];
   assign out_block[28] = inp_block[64-12];
   assign out_block[27] = inp_block[64-52];
   assign out_block[26] = inp_block[64-20];
   assign out_block[25] = inp_block[64-60];   
   assign out_block[24] = inp_block[64-28];   
   assign out_block[23] = inp_block[64-35];
   assign out_block[22] = inp_block[64-3];   
   assign out_block[21] = inp_block[64-43];
   assign out_block[20] = inp_block[64-11];
   assign out_block[19] = inp_block[64-51];
   assign out_block[18] = inp_block[64-19];
   assign out_block[17] = inp_block[64-59];
   assign out_block[16] = inp_block[64-27];   
   assign out_block[15] = inp_block[64-34];
   assign out_block[14] = inp_block[64-2];   
   assign out_block[13] = inp_block[64-42];
   assign out_block[12] = inp_block[64-10];   
   assign out_block[11] = inp_block[64-50];
   assign out_block[10] = inp_block[64-18];
   assign out_block[9] = inp_block[64-58];
   assign out_block[8] = inp_block[64-26];   
   assign out_block[7] = inp_block[64-33];
   assign out_block[6] = inp_block[64-1];
   assign out_block[5] = inp_block[64-41];   
   assign out_block[4] = inp_block[64-9];
   assign out_block[3] = inp_block[64-49];    
   assign out_block[2] = inp_block[64-17];
   assign out_block[1] = inp_block[64-57];
   assign out_block[0] = inp_block[64-25];  

endmodule // FP

module S1_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case ({{inp_bits[5], inp_bits[0]}, inp_bits[4:1]})
	  6'd0  : out_bits = 4'd14;             
	  6'd1  : out_bits = 4'd4;             
	  6'd2  : out_bits = 4'd13;            
	  6'd3  : out_bits = 4'd1;             
	  6'd4  : out_bits = 4'd2;             
	  6'd5  : out_bits = 4'd15;             
	  6'd6  : out_bits = 4'd11;             
	  6'd7  : out_bits = 4'd8;             
	  6'd8  : out_bits = 4'd3;             
	  6'd9  : out_bits = 4'd10;             
	  6'd10 : out_bits = 4'd6;             
	  6'd11 : out_bits = 4'd12;             
	  6'd12 : out_bits = 4'd5;             
	  6'd13 : out_bits = 4'd9;             
	  6'd14 : out_bits = 4'd0;             
	  6'd15 : out_bits = 4'd7;             
	  6'd16 : out_bits = 4'd0;             
	  6'd17 : out_bits = 4'd15;             
	  6'd18 : out_bits = 4'd7;             
	  6'd19 : out_bits = 4'd4;             
	  6'd20 : out_bits = 4'd14;             
	  6'd21 : out_bits = 4'd2;             
	  6'd22 : out_bits = 4'd13;             
	  6'd23 : out_bits = 4'd1;             
	  6'd24 : out_bits = 4'd10;             
	  6'd25 : out_bits = 4'd6;             
	  6'd26 : out_bits = 4'd12;             
	  6'd27 : out_bits = 4'd11;             
	  6'd28 : out_bits = 4'd9;             
	  6'd29 : out_bits = 4'd5;             
	  6'd30 : out_bits = 4'd3;             
	  6'd31 : out_bits = 4'd8;             
	  6'd32 : out_bits = 4'd4;             
	  6'd33 : out_bits = 4'd1;             
	  6'd34 : out_bits = 4'd14;             
	  6'd35 : out_bits = 4'd8;             
	  6'd36 : out_bits = 4'd13;             
	  6'd37 : out_bits = 4'd6;             
	  6'd38 : out_bits = 4'd2;             
	  6'd39 : out_bits = 4'd11;             
	  6'd40 : out_bits = 4'd15;             
	  6'd41 : out_bits = 4'd12;             
	  6'd42 : out_bits = 4'd9;             
	  6'd43 : out_bits = 4'd7;             
	  6'd44 : out_bits = 4'd3;             
	  6'd45 : out_bits = 4'd10;             
	  6'd46 : out_bits = 4'd5;             
	  6'd47 : out_bits = 4'd0;             
	  6'd48 : out_bits = 4'd15;             
	  6'd49 : out_bits = 4'd12;             
	  6'd50 : out_bits = 4'd8;             
	  6'd51 : out_bits = 4'd2;             
	  6'd52 : out_bits = 4'd4;             
	  6'd53 : out_bits = 4'd9;            
	  6'd54 : out_bits = 4'd1;             
	  6'd55 : out_bits = 4'd7;            
	  6'd56 : out_bits = 4'd5;        
	  6'd57 : out_bits = 4'd11;        
	  6'd58 : out_bits = 4'd3;       
	  6'd59 : out_bits = 4'd14;       
	  6'd60 : out_bits = 4'd10;       
	  6'd61 : out_bits = 4'd0;       
	  6'd62 : out_bits = 4'd6;      
	  6'd63 : out_bits = 4'd13;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S1_Box

module S2_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case ({{inp_bits[5], inp_bits[0]}, inp_bits[4:1]})             
	  6'd0  : out_bits = 4'd15;             
	  6'd1  : out_bits = 4'd1;             
	  6'd2  : out_bits = 4'd8;            
	  6'd3  : out_bits = 4'd14;             
	  6'd4  : out_bits = 4'd6;             
	  6'd5  : out_bits = 4'd11;             
	  6'd6  : out_bits = 4'd3;             
	  6'd7  : out_bits = 4'd4;             
	  6'd8  : out_bits = 4'd9;             
	  6'd9  : out_bits = 4'd7;             
	  6'd10 : out_bits = 4'd2;             
	  6'd11 : out_bits = 4'd13;             
	  6'd12 : out_bits = 4'd12;             
	  6'd13 : out_bits = 4'd0;             
	  6'd14 : out_bits = 4'd5;             
	  6'd15 : out_bits = 4'd10;             
	  6'd16 : out_bits = 4'd3;             
	  6'd17 : out_bits = 4'd13;             
	  6'd18 : out_bits = 4'd4;             
	  6'd19 : out_bits = 4'd7;             
	  6'd20 : out_bits = 4'd15;             
	  6'd21 : out_bits = 4'd2;             
	  6'd22 : out_bits = 4'd8;             
	  6'd23 : out_bits = 4'd14;             
	  6'd24 : out_bits = 4'd12;             
	  6'd25 : out_bits = 4'd0;             
	  6'd26 : out_bits = 4'd1;             
	  6'd27 : out_bits = 4'd10;             
	  6'd28 : out_bits = 4'd6;             
	  6'd29 : out_bits = 4'd9;             
	  6'd30 : out_bits = 4'd11;             
	  6'd31 : out_bits = 4'd5;             
	  6'd32 : out_bits = 4'd0;             
	  6'd33 : out_bits = 4'd14;             
	  6'd34 : out_bits = 4'd7;             
	  6'd35 : out_bits = 4'd11;             
	  6'd36 : out_bits = 4'd10;             
	  6'd37 : out_bits = 4'd4;             
	  6'd38 : out_bits = 4'd13;             
	  6'd39 : out_bits = 4'd1;             
	  6'd40 : out_bits = 4'd5;             
	  6'd41 : out_bits = 4'd8;             
	  6'd42 : out_bits = 4'd12;             
	  6'd43 : out_bits = 4'd6;             
	  6'd44 : out_bits = 4'd9;             
	  6'd45 : out_bits = 4'd3;             
	  6'd46 : out_bits = 4'd2;             
	  6'd47 : out_bits = 4'd15;             
	  6'd48 : out_bits = 4'd13;             
	  6'd49 : out_bits = 4'd8;             
	  6'd50 : out_bits = 4'd10;             
	  6'd51 : out_bits = 4'd1;             
	  6'd52 : out_bits = 4'd3;             
	  6'd53 : out_bits = 4'd15;            
	  6'd54 : out_bits = 4'd4;             
	  6'd55 : out_bits = 4'd2;            
	  6'd56 : out_bits = 4'd11;        
	  6'd57 : out_bits = 4'd6;        
	  6'd58 : out_bits = 4'd7;       
	  6'd59 : out_bits = 4'd12;       
	  6'd60 : out_bits = 4'd0;       
	  6'd61 : out_bits = 4'd5;       
	  6'd62 : out_bits = 4'd14;      
	  6'd63 : out_bits = 4'd9;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S2_Box

module S3_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case ({{inp_bits[5], inp_bits[0]}, inp_bits[4:1]})
	  6'd0  : out_bits = 4'd10;             
	  6'd1  : out_bits = 4'd0;             
	  6'd2  : out_bits = 4'd9;            
	  6'd3  : out_bits = 4'd14;             
	  6'd4  : out_bits = 4'd6;             
	  6'd5  : out_bits = 4'd3;             
	  6'd6  : out_bits = 4'd15;             
	  6'd7  : out_bits = 4'd5;             
	  6'd8  : out_bits = 4'd1;             
	  6'd9  : out_bits = 4'd13;             
	  6'd10 : out_bits = 4'd12;             
	  6'd11 : out_bits = 4'd7;             
	  6'd12 : out_bits = 4'd11;             
	  6'd13 : out_bits = 4'd4;             
	  6'd14 : out_bits = 4'd2;             
	  6'd15 : out_bits = 4'd8;             
	  6'd16 : out_bits = 4'd13;             
	  6'd17 : out_bits = 4'd7;             
	  6'd18 : out_bits = 4'd0;             
	  6'd19 : out_bits = 4'd9;             
	  6'd20 : out_bits = 4'd3;             
	  6'd21 : out_bits = 4'd4;             
	  6'd22 : out_bits = 4'd6;             
	  6'd23 : out_bits = 4'd10;             
	  6'd24 : out_bits = 4'd2;             
	  6'd25 : out_bits = 4'd8;             
	  6'd26 : out_bits = 4'd5;             
	  6'd27 : out_bits = 4'd14;             
	  6'd28 : out_bits = 4'd12;             
	  6'd29 : out_bits = 4'd11;             
	  6'd30 : out_bits = 4'd15;             
	  6'd31 : out_bits = 4'd1;             
	  6'd32 : out_bits = 4'd13;             
	  6'd33 : out_bits = 4'd6;             
	  6'd34 : out_bits = 4'd4;             
	  6'd35 : out_bits = 4'd9;             
	  6'd36 : out_bits = 4'd8;             
	  6'd37 : out_bits = 4'd15;             
	  6'd38 : out_bits = 4'd3;             
	  6'd39 : out_bits = 4'd0;             
	  6'd40 : out_bits = 4'd11;             
	  6'd41 : out_bits = 4'd1;             
	  6'd42 : out_bits = 4'd2;             
	  6'd43 : out_bits = 4'd12;             
	  6'd44 : out_bits = 4'd5;             
	  6'd45 : out_bits = 4'd10;             
	  6'd46 : out_bits = 4'd14;             
	  6'd47 : out_bits = 4'd7;             
	  6'd48 : out_bits = 4'd1;             
	  6'd49 : out_bits = 4'd10;             
	  6'd50 : out_bits = 4'd13;             
	  6'd51 : out_bits = 4'd0;             
	  6'd52 : out_bits = 4'd6;             
	  6'd53 : out_bits = 4'd9;            
	  6'd54 : out_bits = 4'd8;             
	  6'd55 : out_bits = 4'd7;            
	  6'd56 : out_bits = 4'd4;        
	  6'd57 : out_bits = 4'd15;        
	  6'd58 : out_bits = 4'd14;       
	  6'd59 : out_bits = 4'd3;       
	  6'd60 : out_bits = 4'd11;       
	  6'd61 : out_bits = 4'd5;       
	  6'd62 : out_bits = 4'd2;      
	  6'd63 : out_bits = 4'd12;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S3_Box

module S4_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case ({{inp_bits[5], inp_bits[0]}, inp_bits[4:1]})   
	  6'd0  : out_bits = 4'd7;             
	  6'd1  : out_bits = 4'd13;             
	  6'd2  : out_bits = 4'd14;            
	  6'd3  : out_bits = 4'd3;             
	  6'd4  : out_bits = 4'd0;             
	  6'd5  : out_bits = 4'd6;             
	  6'd6  : out_bits = 4'd9;             
	  6'd7  : out_bits = 4'd10;             
	  6'd8  : out_bits = 4'd1;             
	  6'd9  : out_bits = 4'd2;             
	  6'd10 : out_bits = 4'd8;             
	  6'd11 : out_bits = 4'd5;             
	  6'd12 : out_bits = 4'd11;             
	  6'd13 : out_bits = 4'd12;             
	  6'd14 : out_bits = 4'd4;             
	  6'd15 : out_bits = 4'd15;             
	  6'd16 : out_bits = 4'd13;             
	  6'd17 : out_bits = 4'd8;             
	  6'd18 : out_bits = 4'd11;             
	  6'd19 : out_bits = 4'd5;             
	  6'd20 : out_bits = 4'd6;             
	  6'd21 : out_bits = 4'd15;             
	  6'd22 : out_bits = 4'd0;             
	  6'd23 : out_bits = 4'd3;             
	  6'd24 : out_bits = 4'd4;             
	  6'd25 : out_bits = 4'd7;             
	  6'd26 : out_bits = 4'd2;             
	  6'd27 : out_bits = 4'd12;             
	  6'd28 : out_bits = 4'd1;             
	  6'd29 : out_bits = 4'd10;             
	  6'd30 : out_bits = 4'd14;             
	  6'd31 : out_bits = 4'd9;             
	  6'd32 : out_bits = 4'd10;             
	  6'd33 : out_bits = 4'd6;             
	  6'd34 : out_bits = 4'd9;             
	  6'd35 : out_bits = 4'd0;             
	  6'd36 : out_bits = 4'd12;             
	  6'd37 : out_bits = 4'd11;             
	  6'd38 : out_bits = 4'd7;             
	  6'd39 : out_bits = 4'd13;             
	  6'd40 : out_bits = 4'd15;             
	  6'd41 : out_bits = 4'd1;             
	  6'd42 : out_bits = 4'd3;             
	  6'd43 : out_bits = 4'd14;             
	  6'd44 : out_bits = 4'd5;             
	  6'd45 : out_bits = 4'd2;             
	  6'd46 : out_bits = 4'd8;             
	  6'd47 : out_bits = 4'd4;             
	  6'd48 : out_bits = 4'd3;             
	  6'd49 : out_bits = 4'd15;             
	  6'd50 : out_bits = 4'd0;             
	  6'd51 : out_bits = 4'd6;             
	  6'd52 : out_bits = 4'd10;             
	  6'd53 : out_bits = 4'd1;            
	  6'd54 : out_bits = 4'd13;             
	  6'd55 : out_bits = 4'd8;            
	  6'd56 : out_bits = 4'd9;        
	  6'd57 : out_bits = 4'd4;        
	  6'd58 : out_bits = 4'd5;       
	  6'd59 : out_bits = 4'd11;       
	  6'd60 : out_bits = 4'd12;       
	  6'd61 : out_bits = 4'd7;       
	  6'd62 : out_bits = 4'd2;      
	  6'd63 : out_bits = 4'd14;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S4_Box

module S5_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case ({{inp_bits[5], inp_bits[0]}, inp_bits[4:1]})   
	  6'd0  : out_bits = 4'd2;             
	  6'd1  : out_bits = 4'd12;             
	  6'd2  : out_bits = 4'd4;            
	  6'd3  : out_bits = 4'd1;             
	  6'd4  : out_bits = 4'd7;             
	  6'd5  : out_bits = 4'd10;             
	  6'd6  : out_bits = 4'd11;             
	  6'd7  : out_bits = 4'd6;             
	  6'd8  : out_bits = 4'd8;             
	  6'd9  : out_bits = 4'd5;             
	  6'd10 : out_bits = 4'd3;             
	  6'd11 : out_bits = 4'd15;             
	  6'd12 : out_bits = 4'd13;             
	  6'd13 : out_bits = 4'd0;             
	  6'd14 : out_bits = 4'd14;             
	  6'd15 : out_bits = 4'd9;             
	  6'd16 : out_bits = 4'd14;             
	  6'd17 : out_bits = 4'd11;             
	  6'd18 : out_bits = 4'd2;             
	  6'd19 : out_bits = 4'd12;             
	  6'd20 : out_bits = 4'd4;             
	  6'd21 : out_bits = 4'd7;             
	  6'd22 : out_bits = 4'd13;             
	  6'd23 : out_bits = 4'd1;             
	  6'd24 : out_bits = 4'd5;             
	  6'd25 : out_bits = 4'd0;             
	  6'd26 : out_bits = 4'd15;             
	  6'd27 : out_bits = 4'd10;             
	  6'd28 : out_bits = 4'd3;             
	  6'd29 : out_bits = 4'd9;             
	  6'd30 : out_bits = 4'd8;             
	  6'd31 : out_bits = 4'd6;             
	  6'd32 : out_bits = 4'd4;             
	  6'd33 : out_bits = 4'd2;             
	  6'd34 : out_bits = 4'd1;             
	  6'd35 : out_bits = 4'd11;             
	  6'd36 : out_bits = 4'd10;             
	  6'd37 : out_bits = 4'd13;             
	  6'd38 : out_bits = 4'd7;             
	  6'd39 : out_bits = 4'd8;             
	  6'd40 : out_bits = 4'd15;             
	  6'd41 : out_bits = 4'd9;             
	  6'd42 : out_bits = 4'd12;             
	  6'd43 : out_bits = 4'd5;             
	  6'd44 : out_bits = 4'd6;             
	  6'd45 : out_bits = 4'd3;             
	  6'd46 : out_bits = 4'd0;             
	  6'd47 : out_bits = 4'd14;             
	  6'd48 : out_bits = 4'd11;             
	  6'd49 : out_bits = 4'd8;             
	  6'd50 : out_bits = 4'd12;             
	  6'd51 : out_bits = 4'd7;             
	  6'd52 : out_bits = 4'd1;             
	  6'd53 : out_bits = 4'd14;            
	  6'd54 : out_bits = 4'd2;             
	  6'd55 : out_bits = 4'd13;            
	  6'd56 : out_bits = 4'd6;        
	  6'd57 : out_bits = 4'd15;        
	  6'd58 : out_bits = 4'd0;       
	  6'd59 : out_bits = 4'd9;       
	  6'd60 : out_bits = 4'd10;       
	  6'd61 : out_bits = 4'd4;       
	  6'd62 : out_bits = 4'd5;      
	  6'd63 : out_bits = 4'd3;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S5_Box

module S6_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case ({{inp_bits[5], inp_bits[0]}, inp_bits[4:1]})   
	  6'd0  : out_bits = 4'd12;             
	  6'd1  : out_bits = 4'd1;             
	  6'd2  : out_bits = 4'd10;            
	  6'd3  : out_bits = 4'd15;             
	  6'd4  : out_bits = 4'd9;             
	  6'd5  : out_bits = 4'd2;             
	  6'd6  : out_bits = 4'd6;             
	  6'd7  : out_bits = 4'd8;             
	  6'd8  : out_bits = 4'd0;             
	  6'd9  : out_bits = 4'd13;             
	  6'd10 : out_bits = 4'd3;             
	  6'd11 : out_bits = 4'd4;             
	  6'd12 : out_bits = 4'd14;             
	  6'd13 : out_bits = 4'd7;             
	  6'd14 : out_bits = 4'd5;             
	  6'd15 : out_bits = 4'd11;             
	  6'd16 : out_bits = 4'd10;             
	  6'd17 : out_bits = 4'd15;             
	  6'd18 : out_bits = 4'd4;             
	  6'd19 : out_bits = 4'd2;             
	  6'd20 : out_bits = 4'd7;             
	  6'd21 : out_bits = 4'd12;             
	  6'd22 : out_bits = 4'd9;             
	  6'd23 : out_bits = 4'd5;             
	  6'd24 : out_bits = 4'd6;             
	  6'd25 : out_bits = 4'd1;             
	  6'd26 : out_bits = 4'd13;             
	  6'd27 : out_bits = 4'd14;             
	  6'd28 : out_bits = 4'd0;             
	  6'd29 : out_bits = 4'd11;             
	  6'd30 : out_bits = 4'd3;             
	  6'd31 : out_bits = 4'd8;             
	  6'd32 : out_bits = 4'd9;             
	  6'd33 : out_bits = 4'd14;             
	  6'd34 : out_bits = 4'd15;             
	  6'd35 : out_bits = 4'd5;             
	  6'd36 : out_bits = 4'd2;             
	  6'd37 : out_bits = 4'd8;             
	  6'd38 : out_bits = 4'd12;             
	  6'd39 : out_bits = 4'd3;             
	  6'd40 : out_bits = 4'd7;             
	  6'd41 : out_bits = 4'd0;             
	  6'd42 : out_bits = 4'd4;             
	  6'd43 : out_bits = 4'd10;             
	  6'd44 : out_bits = 4'd1;             
	  6'd45 : out_bits = 4'd13;             
	  6'd46 : out_bits = 4'd11;             
	  6'd47 : out_bits = 4'd6;             
	  6'd48 : out_bits = 4'd4;             
	  6'd49 : out_bits = 4'd3;             
	  6'd50 : out_bits = 4'd2;             
	  6'd51 : out_bits = 4'd12;             
	  6'd52 : out_bits = 4'd9;             
	  6'd53 : out_bits = 4'd5;            
	  6'd54 : out_bits = 4'd15;             
	  6'd55 : out_bits = 4'd10;            
	  6'd56 : out_bits = 4'd11;        
	  6'd57 : out_bits = 4'd14;        
	  6'd58 : out_bits = 4'd1;       
	  6'd59 : out_bits = 4'd7;       
	  6'd60 : out_bits = 4'd6;       
	  6'd61 : out_bits = 4'd0;       
	  6'd62 : out_bits = 4'd8;      
	  6'd63 : out_bits = 4'd13;	  
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S6_Box

module S7_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case ({{inp_bits[5], inp_bits[0]}, inp_bits[4:1]})   
	  6'd0  : out_bits = 4'd4;             
	  6'd1  : out_bits = 4'd11;             
	  6'd2  : out_bits = 4'd2;            
	  6'd3  : out_bits = 4'd14;             
	  6'd4  : out_bits = 4'd15;             
	  6'd5  : out_bits = 4'd0;             
	  6'd6  : out_bits = 4'd8;             
	  6'd7  : out_bits = 4'd13;             
	  6'd8  : out_bits = 4'd3;             
	  6'd9  : out_bits = 4'd12;             
	  6'd10 : out_bits = 4'd9;             
	  6'd11 : out_bits = 4'd7;             
	  6'd12 : out_bits = 4'd5;             
	  6'd13 : out_bits = 4'd10;             
	  6'd14 : out_bits = 4'd6;             
	  6'd15 : out_bits = 4'd1;             
	  6'd16 : out_bits = 4'd13;             
	  6'd17 : out_bits = 4'd0;             
	  6'd18 : out_bits = 4'd11;             
	  6'd19 : out_bits = 4'd7;             
	  6'd20 : out_bits = 4'd4;             
	  6'd21 : out_bits = 4'd9;             
	  6'd22 : out_bits = 4'd1;             
	  6'd23 : out_bits = 4'd10;             
	  6'd24 : out_bits = 4'd14;             
	  6'd25 : out_bits = 4'd3;             
	  6'd26 : out_bits = 4'd5;             
	  6'd27 : out_bits = 4'd12;             
	  6'd28 : out_bits = 4'd2;             
	  6'd29 : out_bits = 4'd15;             
	  6'd30 : out_bits = 4'd8;             
	  6'd31 : out_bits = 4'd6;             
	  6'd32 : out_bits = 4'd1;             
	  6'd33 : out_bits = 4'd4;             
	  6'd34 : out_bits = 4'd11;             
	  6'd35 : out_bits = 4'd13;             
	  6'd36 : out_bits = 4'd12;             
	  6'd37 : out_bits = 4'd3;             
	  6'd38 : out_bits = 4'd7;             
	  6'd39 : out_bits = 4'd14;             
	  6'd40 : out_bits = 4'd10;             
	  6'd41 : out_bits = 4'd15;             
	  6'd42 : out_bits = 4'd6;             
	  6'd43 : out_bits = 4'd8;             
	  6'd44 : out_bits = 4'd0;             
	  6'd45 : out_bits = 4'd5;             
	  6'd46 : out_bits = 4'd9;             
	  6'd47 : out_bits = 4'd2;             
	  6'd48 : out_bits = 4'd6;             
	  6'd49 : out_bits = 4'd11;             
	  6'd50 : out_bits = 4'd13;             
	  6'd51 : out_bits = 4'd8;             
	  6'd52 : out_bits = 4'd1;             
	  6'd53 : out_bits = 4'd4;            
	  6'd54 : out_bits = 4'd10;             
	  6'd55 : out_bits = 4'd7;            
	  6'd56 : out_bits = 4'd9;        
	  6'd57 : out_bits = 4'd5;        
	  6'd58 : out_bits = 4'd0;       
	  6'd59 : out_bits = 4'd15;       
	  6'd60 : out_bits = 4'd14;       
	  6'd61 : out_bits = 4'd2;       
	  6'd62 : out_bits = 4'd3;      
	  6'd63 : out_bits = 4'd12;  
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S7_Box

module S8_Box (inp_bits, out_bits);

   input logic [5:0] inp_bits;
   output logic [3:0] out_bits;

   always_comb
     begin
	case ({{inp_bits[5], inp_bits[0]}, inp_bits[4:1]})   
	  6'd0  : out_bits = 4'd13;             
	  6'd1  : out_bits = 4'd2;             
	  6'd2  : out_bits = 4'd8;            
	  6'd3  : out_bits = 4'd4;             
	  6'd4  : out_bits = 4'd6;             
	  6'd5  : out_bits = 4'd15;             
	  6'd6  : out_bits = 4'd11;             
	  6'd7  : out_bits = 4'd1;             
	  6'd8  : out_bits = 4'd10;             
	  6'd9  : out_bits = 4'd9;             
	  6'd10 : out_bits = 4'd3;             
	  6'd11 : out_bits = 4'd14;             
	  6'd12 : out_bits = 4'd5;             
	  6'd13 : out_bits = 4'd0;             
	  6'd14 : out_bits = 4'd12;             
	  6'd15 : out_bits = 4'd7;             
	  6'd16 : out_bits = 4'd1;             
	  6'd17 : out_bits = 4'd15;             
	  6'd18 : out_bits = 4'd13;             
	  6'd19 : out_bits = 4'd8;             
	  6'd20 : out_bits = 4'd10;             
	  6'd21 : out_bits = 4'd3;             
	  6'd22 : out_bits = 4'd7;             
	  6'd23 : out_bits = 4'd4;             
	  6'd24 : out_bits = 4'd12;             
	  6'd25 : out_bits = 4'd5;             
	  6'd26 : out_bits = 4'd6;             
	  6'd27 : out_bits = 4'd11;             
	  6'd28 : out_bits = 4'd0;             
	  6'd29 : out_bits = 4'd14;             
	  6'd30 : out_bits = 4'd9;             
	  6'd31 : out_bits = 4'd2;             
	  6'd32 : out_bits = 4'd7;             
	  6'd33 : out_bits = 4'd11;             
	  6'd34 : out_bits = 4'd4;             
	  6'd35 : out_bits = 4'd1;             
	  6'd36 : out_bits = 4'd9;             
	  6'd37 : out_bits = 4'd12;             
	  6'd38 : out_bits = 4'd14;             
	  6'd39 : out_bits = 4'd2;             
	  6'd40 : out_bits = 4'd0;             
	  6'd41 : out_bits = 4'd6;             
	  6'd42 : out_bits = 4'd10;             
	  6'd43 : out_bits = 4'd13;             
	  6'd44 : out_bits = 4'd15;             
	  6'd45 : out_bits = 4'd3;             
	  6'd46 : out_bits = 4'd5;             
	  6'd47 : out_bits = 4'd8;             
	  6'd48 : out_bits = 4'd2;             
	  6'd49 : out_bits = 4'd1;             
	  6'd50 : out_bits = 4'd14;             
	  6'd51 : out_bits = 4'd7;             
	  6'd52 : out_bits = 4'd4;             
	  6'd53 : out_bits = 4'd10;            
	  6'd54 : out_bits = 4'd8;             
	  6'd55 : out_bits = 4'd13;            
	  6'd56 : out_bits = 4'd15;        
	  6'd57 : out_bits = 4'd12;        
	  6'd58 : out_bits = 4'd9;       
	  6'd59 : out_bits = 4'd0;       
	  6'd60 : out_bits = 4'd3;       
	  6'd61 : out_bits = 4'd5;       
	  6'd62 : out_bits = 4'd6;      
	  6'd63 : out_bits = 4'd11;      
	  default : out_bits = 4'd0; 		
        endcase
     end // always_comb
   
endmodule // S8_Box

module DES (input logic [63:0] key, input logic [63:0] plaintext, 
	    input logic encrypt, output logic [63:0] ciphertext);

   logic [47:0] 	SubKey1, SubKey2, SubKey3, SubKey4;   
   logic [47:0] 	SubKey5, SubKey6, SubKey7, SubKey8;   
   logic [47:0] 	SubKey9, SubKey10, SubKey11, SubKey12;
   logic [47:0] 	SubKey13, SubKey14, SubKey15, SubKey16;

<<<<<<< HEAD
   logic [47:0]   sk1, sk2, sk3, sk4;
   logic [47:0]   sk5, sk6, sk7, sk8;
   logic [47:0]   sk9, sk10, sk11, sk12;
   logic [47:0]   sk13, sk14, sk15, sk16;

   logic [63:0]  	ip_out;   
   logic [63:0]   r16_out = 64'h0;   

   logic [63:0]   out1, out2, out3, out4;
   logic [63:0]   out5, out6, out7, out8;
   logic [63:0]   out9, out10, out11, out12;
   logic [63:0]   out13, out14, out15, out16;
=======
   logic [47:0]     sk1, sk2, sk3, sk4;
   logic [47:0]     sk5, sk6, sk7, sk8;
   logic [47:0]     sk9, sk10, sk11, sk12;
   logic [47:0]     sk13, sk14, sk15, sk16;

   logic [63:0] 	ip_out;   
   logic [63:0] 	r16_out = 64'h0;   
>>>>>>> 2cb05479a716221d24a2dce71af84162bc87bae0
   
   // SubKey generation
   GenerateKeys k1 (key, SubKey1, SubKey2, SubKey3, SubKey4,
		    SubKey5, SubKey6, SubKey7, SubKey8,
		    SubKey9, SubKey10, SubKey11, SubKey12,
		    SubKey13, SubKey14, SubKey15, SubKey16);
   // encrypt (encrypt=1) or decrypt (encrypt=0) 
   assign{sk1,sk2,sk3,sk4,sk5,sk6,sk7,sk8,sk9,sk10,sk11,sk12,sk13,sk14,sk15,sk16} = encrpyt ? {SubKey1, SubKey2, SubKey3, SubKey4, SubKey5, SubKey6, SubKey7, SubKey8, SubKey9, SubKey10, SubKey11, SubKey12, SubKey13, SubKey14, SubKey15, SubKey16}:{SubKey16,SubKey15,SubKey14,SubKey13,SubKey12,SubKey11,SubKey10,SubKey9,SubKey8,SubKey7,SubKey6,SubKey5,SubKey4,SubKey3,SubKey2,SubKey1};
   // Initial Permutation (IP)
<<<<<<< HEAD
   IP b1 (plaintext, ip_out); //scrambles
   //round 1
   round r1 (ip_out, sk1, out1); //feistaled block with sk the combined right and left blocks
   // round 2
   round r2 (out1, sk2, out2);
   // round 3
   round r3 (out2, sk3, out3);
   // round 4
   round r4 (out3, sk4, out4);
   // round 5
   round r5 (out4, sk5, out5);
   // round 6
   round r6 (out5, sk6, out6);
   // round 7
   round r7 (out6, sk7, out7);
   // round 8
   round r8 (out7, sk8, out8);
   // round 9
   round r9 (out8, sk9, out9);
   // round 10
   round r10 (out9, sk10, out10);
   // round 11
   round r11 (out10, sk11, out11);
   // round 12
   round r12 (out11, sk12, out12);
   // round 13
   round r13 (out12, sk13, out13);
   // round 14
   round r14 (out13, sk14, out14);
   // round 15
   round r15 (out14, sk15, out15);
   // round 16
   round r16 (out15, sk16, out16);
=======
   IP b1 (plaintext, ip_out);
   // round 1
   logic [63:0] out1;
   round r_1(ip_out, sk1, out1);
   // round 2
   logic [63:0] out2;
   round r_2(out1, sk2, out2);
   // round 3
   logic [63:0] out3;
   round r_3(out2, sk3, out3);
   // round 4
   logic [63:0] out4;
   round r_2(out3, sk4, out4);
   // round 5
   logic [63:0] out5;
   round r_2(out4, sk5, out5);
   // round 6
   logic [63:0] out6;
   round r_2(out5, sk6, out6);
   // round 7
   logic [63:0] out7;
   round r_2(out6, sk7, out7);
   // round 8
   logic [63:0] out8;
   round r_2(out7, sk8, out8);
   // round 9
   logic [63:0] out9;
   round r_2(out8, sk9, out9);
   // round 10
   logic [63:0] out10;
   round r_2(out9, sk10, out10);
   // round 11
   logic [63:0] out11;
   round r_2(out10, sk11, out11);
   // round 12
   logic [63:0] out12;
   round r_2(out11, sk12, out12);
   // round 13
   logic [63:0] out13;
   round r_2(out12, sk13, out13);
   // round 14
   logic [63:0] out14;
   round r_2(out13, sk14, out14);
   // round 15
   logic [63:0] out15;
   round r_2(out14, sk15, out15);
   // round 16
   logic [63:0] out16;
   round r_2(out15, sk16, out16);
>>>>>>> 2cb05479a716221d24a2dce71af84162bc87bae0
   // Final Permutation (IP^{-1}) (swap output of round16)
   FP FP(out16, ciphertext);
   
endmodule // DES